** Profile: "SCHEMATIC1-sim"  [ C:\Users\Amy\Desktop\facultatea masii\Proiect Amelia - V1\proiect amelia - schema reala-PSpiceFiles\SCHEMATIC1\sim.sim ] 

** Creating circuit file "sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/../../Cadence/SPB_17.2/tools/pspice/library/nom.lib" 
.LIB "C:/../../Cadence/SPB_17.2/tools/pspice/library/nomd.lib" 
.LIB "C:/../../Cadence/SPB_17.2/tools/pspice/library/pwrbjt.lib" 
.LIB "C:/../../Cadence/SPB_17.2/tools/pspice/library/phil_diode.lib" 
.LIB "C:/../../Cadence/SPB_17.2/tools/pspice/library/on_bjt.lib" 
.LIB "C:/../../Cadence/SPB_17.2/tools/pspice/library/infineon_s_afbjt.lib" 
.LIB "C:/../../Cadence/SPB_17.2/tools/pspice/library/phil_bjt.lib" 
.LIB "../../../mjd32c.lib" 
.LIB "../../../mjd31c.lib" 
* From [PSPICE NETLIST] section of C:\Users\Amy\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
